module ldpc_encoder_wrapper (
    input           clk,
    input           reset,
    input [359:0]   lpdc_bit_in,
    output [359:0]  lpdc_bit_out
);



endmodule